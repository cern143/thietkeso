module display (start, disable_c, disable_h, mode, clk, rst_n);

input start, disable_c, disable_h, clk, rst_n;

