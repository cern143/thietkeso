module top;

imem  

endmodule
