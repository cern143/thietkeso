module fsm_tb;
